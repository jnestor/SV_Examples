module black(
    input logic pl, pr, gl, gr
    );


endmodule
