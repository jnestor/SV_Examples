//-----------------------------------------------------------------------------
// Module Name   : 
// Project       :
//-----------------------------------------------------------------------------
// Author        :
// Created       :
//-----------------------------------------------------------------------------
// Description   :
//-----------------------------------------------------------------------------
