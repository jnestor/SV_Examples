module black(
    input logic pl, pr, gl, gr
    output logic pc, gc
    );



endmodule
