module black();


endmodule
